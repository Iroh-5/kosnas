component nas.CryptoModule

endpoints {
    CryptoModule: nas.CryptoModule
}
