component nas.CredStorageReader

endpoints {
    CredStorageReader: nas.CredStorageReader
}
