component nas.FsReader

endpoints {
    FsReader: nas.FsReader
}
