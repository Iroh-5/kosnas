component nas.CredStorageWriter

endpoints {
    CredStorageWriter: nas.CredStorageWriter
}
