component nas.FsWriter

endpoints {
    FsWriter: nas.FsWriter
}
